module ALU (
            input [7:0]  A,
            input [7:0]  B,
            input [3:0]  FN,
            output [7:0] result,
            output       overflow,
            output       sign
            );



endmodule
