module seven_segment_driver (
                             input        clk,
                             input        rst_n,
                             input [9:0]  BCD_digit,
                             input        sign,
                             input        overflow,
                             output [3:0] digit_anode,
                             output [6:0] segment
                             );



endmodule
