module synchronizer(
    input clk,
    input reset_n,
    input unsynched,
    output synched
);



endmodule