module binary_to_bcd (
                      input [7:0]  binary_in,
                      output [9:0] bcd_out
                      );



endmodule
