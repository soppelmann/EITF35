module binary_to_sg
  (input  [3:0] binary_in,
   output [7:0] sev_seg);

endmodule
