module keyboard_controller(
    input clk,
    input reset_n,
    input valid_scan_code,
    input [7:0] scan_code,
    output [31:0] scan_codes
);



endmodule
