module debouncer (
                  input  clk,
                  input  rst_n,
                  input  button_in,
                  output button_out
                  );

   reg [19:0] count;
   reg        button_tmp;



endmodule
