module reg_update (
                   input        clk,
                   input        rst_n,
                   input [1:0]  reg_ctrl,
                   output [7:0] A,
                   output [7:0] B
                   );



endmodule
