module serial_to_scancode(
    input clk,
    input reset_n,
    input sample_ready,
    input serial_data,
    output valid_scan_code,
    output [7:0] scan_code
);



endmodule