module falling_edge_detector(
    input clk,
    input reset_n,
    input in,
    output edge_found
);



endmodule