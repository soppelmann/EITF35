module ALU_ctrl (
                 input        clk,
                 input        rst_n,
                 input        enter,
                 input        sign,
                 output [3:0] func,
                 output [1:0] reg_ctrl
                 );



endmodule
