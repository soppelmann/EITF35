module reg_updater (
                   input        clk,
                   input        rst_n,
                   input [1:0]  reg_ctrl,
                   input [7:0]  sw_input,
                   output [7:0] A,
                   output [7:0] B
                   );



endmodule
