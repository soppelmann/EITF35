getz@MBP14.local.3212